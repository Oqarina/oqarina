(***
 * Oqarina
 * Copyright 2021 Carnegie Mellon University.
 *
 * NO WARRANTY. THIS CARNEGIE MELLON UNIVERSITY AND SOFTWARE ENGINEERING
 * INSTITUTE MATERIAL IS FURNISHED ON AN "AS-IS" BASIS. CARNEGIE MELLON
 * UNIVERSITY MAKES NO WARRANTIES OF ANY KIND, EITHER EXPRESSED OR
 * IMPLIED, AS TO ANY MATTER INCLUDING, BUT NOT LIMITED TO, WARRANTY OF
 * FITNESS FOR PURPOSE OR MERCHANTABILITY, EXCLUSIVITY, OR RESULTS
 * OBTAINED FROM USE OF THE MATERIAL. CARNEGIE MELLON UNIVERSITY DOES NOT
 * MAKE ANY WARRANTY OF ANY KIND WITH RESPECT TO FREEDOM FROM PATENT,
 * TRADEMARK, OR COPYRIGHT INFRINGEMENT.
 *
 * Released under a BSD (SEI)-style license, please see license.txt or
 * contact permission@sei.cmu.edu for full terms.
 *
 * [DISTRIBUTION STATEMENT A] This material has been approved for public
 * release and unlimited distribution.  Please see Copyright notice for
 * non-US Government use and distribution.
 *
 * This Software includes and/or makes use of the following Third-Party
 * Software subject to its own license:
 *
 * 1. Coq theorem prover (https://github.com/coq/coq/blob/master/LICENSE)
 * Copyright 2021 INRIA.
 *
 * 2. Coq JSON (https://github.com/liyishuai/coq-json/blob/comrade/LICENSE)
 * Copyright 2021 Yishuai Li.
 *
 * DM21-0762
***)

Require Import Coq.Logic.FunctionalExtensionality.
Require Import Oqarina.core.identifiers.

(*| This module introduces a definition of total maps derived from
Software Fundations. We opted for this design as Coq standard library for FMaps is probably too heavy for our needs.
|*)

Definition total_map (A : Type) := identifier -> A.

Definition t_empty {A : Type} (v : A) : total_map A :=
  (fun _ => v).

Definition t_update {A : Type} (m : total_map A)
                    (x : identifier) (v : A) :=
  fun x' => if identifier_beq x x' then v else m x'.

Notation "'_' '!->' v" := (t_empty v)
  (at level 100, right associativity).

Notation "x '!->' v ';' m" := (t_update m x v)
                              (at level 100, v at next level, right associativity).

Lemma t_apply_empty : forall (A : Type) (x : identifier) (v : A),
  (_ !-> v) x = v.
Proof.
    intros.
    auto.
Qed.

Theorem identifier_eqb_refl : forall s : identifier,
    identifier_beq s s = true.
Proof.
    intros s.
    apply identifier_beq_eq.
    reflexivity.
Qed.

Lemma t_update_eq : forall A (m: total_map A) x v,
  (t_update m x v) x = v.
Proof.
  intros.
  unfold t_update.
  rewrite identifier_eqb_refl.
  reflexivity.
Qed.

Theorem t_update_neq : forall (A : Type) (m : total_map A) x1 x2 v,
  x1 <> x2 ->
  (x1 !-> v ; m) x2 = m x2.
Proof.
    intros.
    unfold t_update.
    rewrite <- identifier_beq_neq in H.
    rewrite H.
    trivial.
  Qed.

Lemma t_update_shadow : forall (A : Type) (m : total_map A) x v1 v2,
  (x !-> v2 ; x !-> v1 ; m) = (x !-> v2 ; m).
Proof.
    intros.
    unfold t_update.

    (* At this stage, we have to prove some equality of functions, this
    can be further simplified using the extensionality axiom. From there, one can simplfiy the goal (remember) and complete the proof.*)
    extensionality x'.
    remember (identifier_beq x x') as eqb.
    induction eqb ; trivial.
Qed.

(* Collection of maps used accross Oqarina *)

Definition list_identifiers_map := total_map (list identifier).

Definition empty_list_identifiers_map : list_identifiers_map :=
    (_ !-> nil).
